magic
tech sky130A
magscale 1 2
timestamp 1653975496
<< error_s >>
rect 560 410 576 426
rect 644 410 660 426
rect 674 410 680 440
rect 544 394 560 410
rect 660 394 680 410
rect 674 324 680 394
rect 536 300 540 324
rect 674 316 684 324
rect 544 300 560 316
rect 660 300 684 316
rect 310 293 368 299
rect 310 259 322 293
rect 560 284 576 300
rect 644 284 660 300
rect 674 280 680 300
rect 560 276 584 280
rect 636 276 660 280
rect 310 253 368 259
rect 710 244 716 476
rect 54 162 112 168
rect 210 162 268 168
rect 54 128 66 162
rect 210 128 222 162
rect 54 122 112 128
rect 210 122 268 128
rect 260 110 300 112
rect 174 89 230 90
rect 174 75 231 89
rect 174 21 210 75
rect 230 21 231 75
rect 174 18 231 21
rect 174 6 230 18
rect 254 6 260 110
rect 264 108 300 110
rect 264 94 330 108
rect 269 90 330 94
rect 272 18 300 78
rect 306 18 330 90
<< nwell >>
rect 230 560 448 562
rect 230 240 710 560
<< nmos >>
rect 230 6 254 90
<< pmos >>
rect 324 340 354 500
<< ndiff >>
rect 174 78 230 90
rect 174 18 186 78
rect 220 18 230 78
rect 174 6 230 18
rect 254 78 312 90
rect 254 18 266 78
rect 300 18 312 78
rect 254 6 312 18
<< pdiff >>
rect 266 488 324 500
rect 266 352 278 488
rect 312 352 324 488
rect 266 340 324 352
rect 354 488 412 500
rect 354 352 366 488
rect 400 352 412 488
rect 354 340 412 352
<< ndiffc >>
rect 186 18 220 78
rect 266 18 299 78
<< pdiffc >>
rect 278 352 312 488
rect 366 352 400 488
<< psubdiff >>
rect 486 -130 510 -10
rect 660 -130 684 -10
<< nsubdiff >>
rect 540 410 680 440
rect 540 300 560 410
rect 660 300 680 410
rect 540 280 680 300
<< psubdiffcont >>
rect 510 -130 660 -10
<< nsubdiffcont >>
rect 560 300 660 410
<< poly >>
rect 324 500 354 526
rect 50 150 120 310
rect 324 309 354 340
rect 306 293 372 309
rect 306 259 322 293
rect 356 259 372 293
rect 306 243 372 259
rect 310 180 370 243
rect 260 178 370 180
rect 206 162 370 178
rect 206 128 222 162
rect 256 128 370 162
rect 206 112 370 128
rect 224 90 254 112
rect 260 110 370 112
rect 224 -20 254 6
<< polycont >>
rect 322 259 356 293
rect 222 128 256 162
<< locali >>
rect 370 504 420 630
rect 30 500 100 504
rect 278 500 312 504
rect -220 420 100 500
rect 170 488 312 500
rect 170 430 278 488
rect -220 -150 -130 420
rect 278 336 312 352
rect 366 488 420 504
rect 400 440 420 488
rect 366 336 400 352
rect 306 259 322 293
rect 356 259 372 293
rect 206 128 222 162
rect 256 128 272 162
rect 10 10 60 90
rect 186 78 220 94
rect 264 78 308 94
rect 110 18 186 40
rect 299 18 308 78
rect 16 -40 56 10
rect 110 0 220 18
rect 140 -150 180 0
rect 264 -40 308 18
rect 494 -130 510 -10
rect 660 -130 676 -10
rect -220 -210 180 -150
<< viali >>
rect 260 630 440 810
rect 278 352 312 488
rect 366 352 400 488
rect 322 259 356 293
rect 222 128 256 162
rect 186 18 220 78
rect 266 18 299 78
rect 10 -100 70 -40
rect 240 -100 310 -40
<< metal1 >>
rect 248 810 452 816
rect -210 630 260 810
rect 440 630 452 810
rect 248 624 452 630
rect 272 488 318 500
rect 272 352 278 488
rect 312 352 318 488
rect 272 340 318 352
rect 360 488 406 500
rect 360 352 366 488
rect 400 352 406 488
rect 360 340 406 352
rect 310 293 368 299
rect 310 259 322 293
rect 356 259 368 293
rect 310 253 368 259
rect 210 162 268 168
rect 210 128 222 162
rect 256 128 268 162
rect 210 122 268 128
rect 180 78 226 90
rect 180 18 186 78
rect 220 18 226 78
rect 180 6 226 18
rect 260 78 306 90
rect 260 18 266 78
rect 300 18 306 78
rect 260 6 306 18
rect -2 -40 82 -34
rect 228 -40 322 -34
rect -2 -100 10 -40
rect 70 -100 240 -40
rect -2 -106 82 -100
rect 228 -106 240 -100
rect 230 -120 240 -106
rect 310 -106 322 -40
rect 310 -120 320 -106
<< via1 >>
rect 260 630 440 810
rect 10 -100 70 -40
rect 240 -100 310 -40
rect 240 -120 310 -100
<< metal2 >>
rect 260 810 440 820
rect 260 620 440 630
rect 10 -40 70 -30
rect 10 -110 70 -100
rect 240 -40 310 -30
rect 240 -130 310 -120
use sky130_fd_pr__nfet_01v8_A64BNL  sky130_fd_pr__nfet_01v8_A64BNL_0
timestamp 0
transform 1 0 83 0 1 79
box -73 -99 73 99
use sky130_fd_pr__pfet_01v8_L3EZX8  sky130_fd_pr__pfet_01v8_L3EZX8_0
timestamp 1653938479
transform 1 0 139 0 1 384
box -109 -144 109 178
<< labels >>
rlabel metal1 -210 710 -210 710 1 vdd
port 3 n
rlabel poly 50 200 50 200 7 A
port 1 w
rlabel poly 310 220 310 220 7 B
port 2 w
rlabel locali -130 110 -130 110 3 y
port 4 e
rlabel metal1 90 -40 90 -40 5 GND
port 5 s
<< end >>
