**.subckt delay_singlestage
**.ends
** flattened .save nodes
.end
