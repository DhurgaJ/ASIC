magic
tech sky130A
magscale 1 2
timestamp 1653977800
<< error_p >>
rect -109 -144 109 178
<< nwell >>
rect -109 -144 109 178
<< pmos >>
rect -15 -44 15 116
<< pdiff >>
rect -73 104 -15 116
rect -73 -32 -61 104
rect -27 -32 -15 104
rect -73 -44 -15 -32
rect 15 104 73 116
rect 15 -32 27 104
rect 61 -32 73 104
rect 15 -44 73 -32
<< pdiffc >>
rect -61 -32 -27 104
rect 27 -32 61 104
<< poly >>
rect -15 116 15 142
rect -15 -75 15 -44
rect -33 -91 33 -75
rect -33 -125 -17 -91
rect 17 -125 33 -91
rect -33 -141 33 -125
<< polycont >>
rect -17 -125 17 -91
<< locali >>
rect -61 104 -27 120
rect -61 -48 -27 -32
rect 27 104 61 120
rect 27 -48 61 -32
rect -33 -125 -17 -91
rect 17 -125 33 -91
<< viali >>
rect -61 -32 -27 104
rect 27 -32 61 104
rect -17 -125 17 -91
<< metal1 >>
rect -67 104 -21 116
rect -67 -32 -61 104
rect -27 -32 -21 104
rect -67 -44 -21 -32
rect 21 104 67 116
rect 21 -32 27 104
rect 61 -32 67 104
rect 21 -44 67 -32
rect -29 -91 29 -85
rect -29 -125 -17 -91
rect 17 -125 29 -91
rect -29 -131 29 -125
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 0.8 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
